//----------------------------------------------------------------------------
//File Name    : xxx 
//Author       : xxx 
//----------------------------------------------------------------------------
//Module Hierarchy :
//xxx_inst |-xxx
//----------------------------------------------------------------------------
//Release History :
//Version         Date           Author        Description
// 1.0          2019-01-01       xxx			1st draft
//----------------------------------------------------------------------------
//Main Function:
//a)xxx
//b)xxx
//c)xxx
//----------------------------------------------------------------------------
module xxx();

////////////////////////////////////////////////////////////////////////////////////////////////////
//                                                                                                //
//    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __//
// __|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |/
//                                                                                                //
//                                                                                                //
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//		xxx_name																				  //	
////////////////////////////////////////////////////////////////////////////////////////////////////

mkdir -p ~/.vim/template

cp -rf template.v ~/.vim/template.v

sudo gvim /etc/vim/vimrc

autocmd BufNewFile *.v 0r /home/cqiu/.vim/template/template.v

endmodule

