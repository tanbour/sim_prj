//=========================== ZTE Corporation=================================//
//   Information contained in this Confidential and Proprietary work has        
//   been obtained by ZTE Corporation. This Design may be used only as          
//   authorized by a Licensing Agreement from ZTE Corporation.                  
//                                                                              
//            COPYRIGHT (C) 2008 ZTE CORPORATION                                
//                  ALL RIGHTS RESERVED                                         
//                                                                              
//   The entire notice above must be displayed on all authorized ZTE            
//   copies.  Copies may be made only to the extended consent by a              
//   Licensing Agreement from ZTE Corporation.                                  
//----------------------------------------------------------------------------//
//      Project and Control Information	                                       
//----------------------------------------------------------------------------//
//      Project Name              :   crc32_d32                             
//      Last Version              :   2.0                                       
//      This Version              :   2.0                                       
//      This module name          :   crc32_d32.v                           
//      This File generated by    :                                             
//      This File updated by      :   None                                      
//      Updated detail            :   None                                      
//----------------------------------------------------------------------------//
//      ZTE Basic Module(s) Information                                         
//----------------------------------------------------------------------------//
//      Included Contents in this Module                                        
//      File Format                :   Verilog HDL                              
//      Included File Name(s)      :   None                                     
//      Included Module(s) Name    :   None                                     
//      Function Block(s)  Name    :   None                                     
//      Task Block(s) Name         :   None                                     
//----------------------------------------------------------------------------//
//       Overview                                                               
//----------------------------------------------------------------------------//
//    CRC calculation
//      Options:
//        Data Width    : 32
//        CRC Init      : All "1"
//        Byte Reverse  : Enable
//        CRC Level     : 32
//        Polynomial    : x32+x26+x23+x22+x16+x12+x11+x10+x8+x7+x5+x4+x2+x+1
//                        1_0000_0100_1100_0001_0001_1101_1011_0111 [32 -> 0]
//                        CRC-32
//----------------------------------------------------------------------------//

module crc32_d32 (
   c,
   crc_out,
   d,
   calc,
   init,
   d_valid,
   clk,
   reset
   );

input         clk;
input         reset;
input  [31:0]  d;
input         calc;
input         init;
input         d_valid;
output [31:0] c;
output [31:0]  crc_out;

reg    [31:0] c;
reg    [31:0]  crc_out;
wire   [31:0] crc_next;

always @ (posedge clk or posedge reset)
begin
   if (reset) begin
      c <= 32'hFFFFFFFF;
      crc_out <=  32'hFFFFFFFF;
   end
   else if (init) begin
      c <= 32'hFFFFFFFF;
      crc_out <=  32'hFFFFFFFF;
   end
   else if (calc & d_valid) begin
      c <= crc_next;
      crc_out <= ~{crc_next[24], crc_next[25], crc_next[26], crc_next[27], crc_next[28], crc_next[29], crc_next[30], crc_next[31], crc_next[16], crc_next[17], crc_next[18], crc_next[19], crc_next[20], crc_next[21], crc_next[22], crc_next[23], crc_next[8], crc_next[9], crc_next[10], crc_next[11], crc_next[12], crc_next[13], crc_next[14], crc_next[15], crc_next[0], crc_next[1], crc_next[2], crc_next[3], crc_next[4], crc_next[5], crc_next[6], crc_next[7]};
   end
end

  assign crc_next[0] = c[0]^c[6]^c[9]^c[10]^c[12]^c[16]^c[24]^c[25]^c[26]^c[28]^c[29]^c[30]^c[31]^d[1]^d[7]^d[11]^d[13]^d[14]^d[23]^d[24]^d[25]^d[26]^d[27]^d[29]^d[30]^d[31];
  assign crc_next[1] = c[0]^c[1]^c[6]^c[7]^c[9]^c[11]^c[12]^c[13]^c[16]^c[17]^c[24]^c[27]^c[28]^d[0]^d[1]^d[6]^d[7]^d[10]^d[11]^d[12]^d[14]^d[22]^d[23]^d[27]^d[28]^d[31];
  assign crc_next[2] = c[0]^c[1]^c[2]^c[6]^c[7]^c[8]^c[9]^c[13]^c[14]^c[16]^c[17]^c[18]^c[24]^c[26]^c[30]^c[31]^d[0]^d[1]^d[5]^d[6]^d[7]^d[9]^d[10]^d[14]^d[15]^d[21]^d[22]^d[23]^d[24]^d[25]^d[29]^d[31];
  assign crc_next[3] = c[1]^c[2]^c[3]^c[7]^c[8]^c[9]^c[10]^c[14]^c[15]^c[17]^c[18]^c[19]^c[25]^c[27]^c[31]^d[0]^d[4]^d[5]^d[6]^d[8]^d[9]^d[13]^d[14]^d[15]^d[20]^d[21]^d[22]^d[24]^d[28]^d[30];
  assign crc_next[4] = c[0]^c[2]^c[3]^c[4]^c[6]^c[8]^c[11]^c[12]^c[15]^c[18]^c[19]^c[20]^c[24]^c[25]^c[29]^c[30]^c[31]^d[1]^d[3]^d[4]^d[5]^d[7]^d[8]^d[11]^d[12]^d[15]^d[19]^d[20]^d[21]^d[24]^d[25]^d[26]^d[30]^d[31];
  assign crc_next[5] = c[0]^c[1]^c[3]^c[4]^c[5]^c[6]^c[7]^c[10]^c[13]^c[19]^c[20]^c[21]^c[24]^c[28]^c[29]^d[0]^d[1]^d[2]^d[3]^d[4]^d[6]^d[7]^d[10]^d[13]^d[18]^d[19]^d[20]^d[26]^d[27]^d[31];
  assign crc_next[6] = c[1]^c[2]^c[4]^c[5]^c[6]^c[7]^c[8]^c[11]^c[14]^c[20]^c[21]^c[22]^c[25]^c[29]^c[30]^d[0]^d[1]^d[2]^d[3]^d[5]^d[6]^d[9]^d[12]^d[15]^d[17]^d[18]^d[19]^d[25]^d[26]^d[30];
  assign crc_next[7] = c[0]^c[2]^c[3]^c[5]^c[7]^c[8]^c[10]^c[15]^c[16]^c[21]^c[22]^c[23]^c[24]^c[25]^c[28]^c[29]^d[0]^d[2]^d[4]^d[5]^d[7]^d[8]^d[13]^d[15]^d[16]^d[17]^d[18]^d[23]^d[26]^d[27]^d[30]^d[31];
  assign crc_next[8] = c[0]^c[1]^c[3]^c[4]^c[8]^c[10]^c[11]^c[12]^c[17]^c[22]^c[23]^c[28]^c[31]^d[3]^d[4]^d[6]^d[7]^d[11]^d[12]^d[13]^d[15]^d[16]^d[17]^d[22]^d[24]^d[27];
  assign crc_next[9] = c[1]^c[2]^c[4]^c[5]^c[9]^c[11]^c[12]^c[13]^c[18]^c[23]^c[24]^c[29]^d[2]^d[3]^d[5]^d[6]^d[10]^d[11]^d[12]^d[14]^d[16]^d[21]^d[26]^d[31];
  assign crc_next[10] = c[0]^c[2]^c[3]^c[5]^c[9]^c[13]^c[14]^c[16]^c[19]^c[26]^c[28]^c[29]^c[31]^d[2]^d[4]^d[5]^d[7]^d[9]^d[10]^d[14]^d[20]^d[23]^d[24]^d[26]^d[27]^d[29];
  assign crc_next[11] = c[0]^c[1]^c[3]^c[4]^c[9]^c[12]^c[14]^c[15]^c[16]^c[17]^c[20]^c[24]^c[25]^c[26]^c[27]^c[28]^c[31]^d[3]^d[4]^d[6]^d[7]^d[8]^d[9]^d[11]^d[14]^d[19]^d[22]^d[23]^d[24]^d[27]^d[28]^d[29]^d[30]^d[31];
  assign crc_next[12] = c[0]^c[1]^c[2]^c[4]^c[5]^c[6]^c[9]^c[12]^c[13]^c[15]^c[17]^c[18]^c[21]^c[24]^c[27]^c[30]^c[31]^d[1]^d[2]^d[3]^d[5]^d[6]^d[7]^d[8]^d[10]^d[11]^d[14]^d[18]^d[21]^d[22]^d[24]^d[25]^d[28]^d[31];
  assign crc_next[13] = c[1]^c[2]^c[3]^c[5]^c[6]^c[7]^c[10]^c[13]^c[14]^c[16]^c[18]^c[19]^c[22]^c[25]^c[28]^c[31]^d[0]^d[1]^d[2]^d[4]^d[5]^d[6]^d[9]^d[10]^d[13]^d[17]^d[20]^d[21]^d[23]^d[24]^d[27]^d[30];
  assign crc_next[14] = c[2]^c[3]^c[4]^c[6]^c[7]^c[8]^c[11]^c[14]^c[15]^c[17]^c[19]^c[20]^c[23]^c[26]^c[29]^d[0]^d[1]^d[3]^d[4]^d[5]^d[8]^d[9]^d[12]^d[15]^d[16]^d[19]^d[20]^d[22]^d[26]^d[29];
  assign crc_next[15] = c[3]^c[4]^c[5]^c[7]^c[8]^c[9]^c[12]^c[15]^c[16]^c[18]^c[20]^c[21]^c[24]^c[27]^c[30]^d[0]^d[2]^d[3]^d[4]^d[8]^d[11]^d[14]^d[15]^d[18]^d[19]^d[21]^d[23]^d[25]^d[28]^d[31];
  assign crc_next[16] = c[0]^c[4]^c[5]^c[8]^c[12]^c[13]^c[17]^c[19]^c[21]^c[22]^c[24]^c[26]^c[29]^c[30]^d[2]^d[3]^d[7]^d[10]^d[11]^d[15]^d[17]^d[18]^d[20]^d[22]^d[25]^d[26]^d[29]^d[31];
  assign crc_next[17] = c[1]^c[5]^c[6]^c[9]^c[13]^c[14]^c[18]^c[20]^c[22]^c[23]^c[25]^c[27]^c[30]^c[31]^d[1]^d[2]^d[6]^d[9]^d[10]^d[14]^d[16]^d[17]^d[19]^d[21]^d[24]^d[25]^d[28]^d[30];
  assign crc_next[18] = c[2]^c[6]^c[7]^c[10]^c[14]^c[15]^c[19]^c[21]^c[23]^c[24]^c[26]^c[28]^c[31]^d[0]^d[1]^d[5]^d[8]^d[9]^d[13]^d[16]^d[18]^d[20]^d[24]^d[27]^d[29]^d[31];
  assign crc_next[19] = c[3]^c[7]^c[8]^c[11]^c[15]^c[16]^c[20]^c[22]^c[24]^c[25]^c[27]^c[29]^d[0]^d[4]^d[8]^d[12]^d[15]^d[17]^d[19]^d[23]^d[26]^d[28]^d[30]^d[31];
  assign crc_next[20] = c[4]^c[8]^c[9]^c[12]^c[16]^c[17]^c[21]^c[23]^c[25]^c[26]^c[28]^c[30]^d[3]^d[11]^d[14]^d[15]^d[16]^d[18]^d[22]^d[23]^d[25]^d[27]^d[29]^d[30];
  assign crc_next[21] = c[5]^c[9]^c[10]^c[13]^c[17]^c[18]^c[22]^c[24]^c[26]^c[27]^c[29]^c[31]^d[2]^d[10]^d[13]^d[14]^d[17]^d[21]^d[22]^d[24]^d[26]^d[28]^d[29]^d[31];
  assign crc_next[22] = c[0]^c[9]^c[11]^c[12]^c[14]^c[16]^c[18]^c[19]^c[23]^c[24]^c[26]^c[27]^c[29]^c[31]^d[7]^d[9]^d[11]^d[12]^d[14]^d[16]^d[20]^d[21]^d[23]^d[24]^d[26]^d[28]^d[29]^d[31];
  assign crc_next[23] = c[0]^c[1]^c[6]^c[9]^c[13]^c[15]^c[16]^c[17]^c[19]^c[20]^c[26]^c[27]^c[29]^c[31]^d[1]^d[6]^d[7]^d[8]^d[10]^d[14]^d[19]^d[20]^d[22]^d[23]^d[24]^d[26]^d[28]^d[29];
  assign crc_next[24] = c[1]^c[2]^c[7]^c[10]^c[14]^c[16]^c[17]^c[18]^c[20]^c[21]^c[27]^c[28]^c[30]^d[0]^d[5]^d[6]^d[9]^d[13]^d[18]^d[19]^d[21]^d[22]^d[23]^d[25]^d[27]^d[28];
  assign crc_next[25] = c[2]^c[3]^c[8]^c[11]^c[15]^c[17]^c[18]^c[19]^c[21]^c[22]^c[28]^c[29]^c[31]^d[4]^d[5]^d[8]^d[12]^d[15]^d[17]^d[18]^d[20]^d[21]^d[22]^d[24]^d[26]^d[27];
  assign crc_next[26] = c[0]^c[3]^c[4]^c[6]^c[10]^c[18]^c[19]^c[20]^c[22]^c[23]^c[24]^c[25]^c[26]^c[28]^c[31]^d[1]^d[3]^d[4]^d[7]^d[13]^d[16]^d[17]^d[19]^d[20]^d[21]^d[24]^d[27]^d[29]^d[30]^d[31];
  assign crc_next[27] = c[1]^c[4]^c[5]^c[7]^c[11]^c[19]^c[20]^c[21]^c[23]^c[24]^c[25]^c[26]^c[27]^c[29]^d[0]^d[2]^d[3]^d[6]^d[12]^d[16]^d[18]^d[19]^d[20]^d[26]^d[28]^d[29]^d[30]^d[31];
  assign crc_next[28] = c[2]^c[5]^c[6]^c[8]^c[12]^c[20]^c[21]^c[22]^c[24]^c[25]^c[26]^c[27]^c[28]^c[30]^d[1]^d[2]^d[5]^d[11]^d[15]^d[17]^d[18]^d[19]^d[25]^d[27]^d[28]^d[29]^d[30]^d[31];
  assign crc_next[29] = c[3]^c[6]^c[7]^c[9]^c[13]^c[21]^c[22]^c[23]^c[25]^c[26]^c[27]^c[28]^c[29]^c[31]^d[0]^d[1]^d[4]^d[10]^d[14]^d[16]^d[17]^d[18]^d[24]^d[26]^d[27]^d[28]^d[29]^d[30];
  assign crc_next[30] = c[4]^c[7]^c[8]^c[10]^c[14]^c[22]^c[23]^c[24]^c[26]^c[27]^c[28]^c[29]^c[30]^d[0]^d[3]^d[9]^d[13]^d[15]^d[16]^d[17]^d[25]^d[26]^d[27]^d[28]^d[29]^d[31];
  assign crc_next[31] = c[5]^c[8]^c[9]^c[11]^c[15]^c[23]^c[24]^c[25]^c[27]^c[28]^c[29]^c[30]^c[31]^d[2]^d[8]^d[12]^d[14]^d[15]^d[16]^d[24]^d[25]^d[26]^d[27]^d[28]^d[30]^d[31];

endmodule
