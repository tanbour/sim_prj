//--------------------------------------------------------------------------------------------------
//File Name    : sync_clka2clkb 
//Author       : sync_clka2clkb 
//--------------------------------------------------------------------------------------------------
//Module Hierarchy :
//sync_clka2clkb_inst |-sync_clka2clkb
//--------------------------------------------------------------------------------------------------
//Release History :
//Version         Date           Author        		Description
// 1.0          2019-01-01       sync_clka2clkb		1st draft
//--------------------------------------------------------------------------------------------------
//Main Function Tree:
//a)sync_clka2clkb: 
//Description Function:
//sync_clka2clkb
//--------------------------------------------------------------------------------------------------
module sync_clka2clkb();
////////////////////////////////////////////////////////////////////////////////////////////////////
// Naming specification																			  // 
// (1) 											  												  // 
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//                                                                                                //
//    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __//
// __|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |/
//                                                                                                //
//                                                                                                //
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//		sync_clka2clkb_name																		  //	
////////////////////////////////////////////////////////////////////////////////////////////////////

endmodule


