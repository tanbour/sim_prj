//--------------------------------------------------------------------------------------------------
//File Name    : wptr_full 
//Author       : wptr_full 
//--------------------------------------------------------------------------------------------------
//Module Hierarchy :
//wptr_full_inst |-wptr_full
//--------------------------------------------------------------------------------------------------
//Release History :
//Version         Date           Author        Description
// 1.0          2019-01-01       wptr_full			1st draft
//--------------------------------------------------------------------------------------------------
//Main Function Tree:
//a)wptr_full: 
//Description Function:
//wptr_full
//--------------------------------------------------------------------------------------------------
module wptr_full();
////////////////////////////////////////////////////////////////////////////////////////////////////
// Naming specification																			  // 
// (1) 											  												  // 
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//                                                                                                //
//    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __//
// __|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |/
//                                                                                                //
//                                                                                                //
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//		wptr_full_name																			  //	
////////////////////////////////////////////////////////////////////////////////////////////////////

endmodule


