//--------------------------------------------------------------------------------------------------
//File Name    : fifomem 
//Author       : fifomem 
//--------------------------------------------------------------------------------------------------
//Module Hierarchy :
//fifomem_inst |-fifomem
//--------------------------------------------------------------------------------------------------
//Release History :
//Version         Date           Author        Description
// 1.0          2019-01-01       fifomem			1st draft
//--------------------------------------------------------------------------------------------------
//Main Function Tree:
//a)fifomem: 
//Description Function:
//fifomem
//--------------------------------------------------------------------------------------------------
module fifomem();
////////////////////////////////////////////////////////////////////////////////////////////////////
// Naming specification																			  // 
// (1) 											  												  // 
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//                                                                                                //
//    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __//
// __|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |/
//                                                                                                //
//                                                                                                //
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//		fifomem_name																				  //	
////////////////////////////////////////////////////////////////////////////////////////////////////

endmodule


