//--------------------------------------------------------------------------------------------------
//File Name    : rptr_empty 
//Author       : rptr_empty 
//--------------------------------------------------------------------------------------------------
//Module Hierarchy :
//rptr_empty_inst |-rptr_empty
//--------------------------------------------------------------------------------------------------
//Release History :
//Version         Date           Author        Description
// 1.0          2019-01-01       rptr_empty			1st draft
//--------------------------------------------------------------------------------------------------
//Main Function Tree:
//a)rptr_empty: 
//Description Function:
//rptr_empty
//--------------------------------------------------------------------------------------------------
module rptr_empty();
////////////////////////////////////////////////////////////////////////////////////////////////////
// Naming specification																			  // 
// (1) 											  												  // 
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//                                                                                                //
//    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __//
// __|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |/
//                                                                                                //
//                                                                                                //
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//		rptr_empty_name																				  //	
////////////////////////////////////////////////////////////////////////////////////////////////////

endmodule


